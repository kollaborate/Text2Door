https://www.google.com/accounts/ClientLogin - OK
Logged in to Google - Auth token received
https://www.google.com/voice/b/0/settings/tab/phones - OK
https://www.google.com/voice/b/0 - OK
Successfully Received rnr_se.
https://www.google.com/voice/b/0/inbox/recent/sms/unread/ - OK
https://www.google.com/voice/b/0/inbox/recent/sms/unread/ - OK
https://www.google.com/voice/b/0/inbox/recent/sms/unread/ - OK
https://www.google.com/voice/b/0/inbox/recent/sms/unread/ - OK
https://www.google.com/voice/b/0/inbox/recent/sms/unread/ - OK
